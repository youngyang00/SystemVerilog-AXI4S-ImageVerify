`ifndef AXI4S_INTERFACE
`define AXI4S_INTERFACE
interface axi4s_io(input bit clock);
   logic                i_rstn;
   logic [95:0]         s_axis_tdata;
   logic                s_axis_tvalid;
   logic                s_axis_tready;
   logic [95:0]         m_axis_tdata;
   logic                m_axis_tvalid;
   logic                m_axis_tready;
   logic                eol;
   logic                eof;

   clocking cb @(posedge clock);
      default input  #2ns  output #2ns;
      output i_rstn;
      output s_axis_tdata;
      input  s_axis_tready;
      input  m_axis_tdata;
      input  m_axis_tvalid;
      input  eol;
      input  eof;
   endclocking


   clocking signal_drv @(posedge clock);
      default input  #2ns  output #2ns;
      output m_axis_tready;
      output s_axis_tvalid;
   endclocking


   clocking signal_smp @(posedge clock);
      default input  #2ns  output #2ns;
      input m_axis_tready;
      input s_axis_tvalid;
   endclocking

   modport TB (
      clocking cb,
      clocking signal_drv,
      clocking signal_smp
   );
endinterface
`endif
